/***********************************************************************
   cpu datapath
 ***********************************************************************/

